
module IMPOR ( out, out_valid, ready, in, mode, in_valid, clk, rst_n );
  output [2:0] out;
  input [2:0] in;
  input [2:0] mode;
  input in_valid, clk, rst_n;
  output out_valid, ready;
  wire   rst, sta, N53, N54, N55, N58, N59, N60, N61, N62, N63, N64, N65, N67,
         N68, N69, N70, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N91, N92, N93, N94, N95, N404, N405, N406, N419,
         N420, N421, N433, N434, N435, N448, N449, N450, N461, N462, N463,
         N467, N468, N469, N473, N474, N475, N479, N480, N481, n44, n45, n46,
         n47, n49, n50, n51, n52, n53, n54, n55, n56, n57, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, add_x_41_1_carry_2_,
         add_x_41_1_carry_3_, add_x_41_1_carry_4_, add_x_41_1_carry_5_,
         add_x_41_1_carry_6_, add_x_41_1_carry_7_, add_x_41_1_carry_8_,
         add_x_41_1_carry_9_, add_x_41_1_carry_10_, add_x_41_1_carry_11_,
         add_x_41_1_carry_12_, add_x_41_1_carry_14_, add_x_41_1_carry_15_,
         add_x_41_1_carry_16_, add_x_41_1_carry_17_, add_x_41_1_carry_18_,
         add_x_41_1_carry_19_, add_x_41_1_carry_20_, add_x_41_0_carry_2_,
         add_x_41_0_carry_3_, add_x_41_0_carry_6_, add_x_41_0_carry_7_,
         add_x_41_0_carry_8_, add_x_41_0_carry_9_, add_x_41_0_carry_10_,
         add_x_41_0_carry_11_, add_x_41_0_carry_12_, add_x_41_0_carry_13_,
         add_x_41_0_carry_15_, add_x_41_0_carry_16_, add_x_41_0_carry_17_,
         add_x_41_0_carry_18_, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n394, n434, n435;
  wire   [2:0] sta20;
  wire   [2:0] sta21;
  wire   [2:0] sta22;
  wire   [2:0] sta23;
  wire   [2:0] sta24;
  wire   [2:0] sta25;
  wire   [2:0] sta26;
  wire   [2:0] sta27;
  wire   [2:0] sta28;
  wire   [20:0] cnt2;
  wire   [20:0] cnt1;

  OAI21XL U32 ( .A0(n95), .A1(n97), .B0(n105), .Y(n106) );
  OAI22XL U33 ( .A0(mode[2]), .A1(n97), .B0(n95), .B1(mode[1]), .Y(n107) );
  AOI2BB1X1 U35 ( .A0N(n108), .A1N(n97), .B0(n104), .Y(n109) );
  OAI22XL U36 ( .A0(mode[0]), .A1(n83), .B0(n97), .B1(n71), .Y(n110) );
  OAI22XL U38 ( .A0(mode[0]), .A1(n84), .B0(n97), .B1(n72), .Y(n112) );
  OAI22XL U39 ( .A0(mode[0]), .A1(n85), .B0(n97), .B1(n73), .Y(n113) );
  OAI22XL U40 ( .A0(mode[2]), .A1(mode[1]), .B0(n95), .B1(n97), .Y(n114) );
  AOI222XL U50 ( .A0(n113), .A1(n96), .B0(n99), .B1(sta27[0]), .C0(n111), .C1(
        N448), .Y(n121) );
  OAI22XL U51 ( .A0(n109), .A1(n121), .B0(n89), .B1(n79), .Y(N473) );
  AOI222XL U52 ( .A0(n112), .A1(n96), .B0(n99), .B1(sta27[1]), .C0(n111), .C1(
        N449), .Y(n122) );
  OAI22XL U53 ( .A0(n109), .A1(n122), .B0(n89), .B1(n78), .Y(N474) );
  AOI222XL U54 ( .A0(n110), .A1(n96), .B0(n99), .B1(sta27[2]), .C0(n111), .C1(
        N450), .Y(n123) );
  OAI22XL U55 ( .A0(n109), .A1(n123), .B0(n89), .B1(n77), .Y(N475) );
  AOI222XL U56 ( .A0(n99), .A1(sta21[0]), .B0(n90), .B1(sta25[0]), .C0(n108), 
        .C1(N404), .Y(n124) );
  OAI222XL U57 ( .A0(n64), .A1(n88), .B0(n73), .B1(n107), .C0(n97), .C1(n124), 
        .Y(N467) );
  AOI222XL U58 ( .A0(n99), .A1(sta21[1]), .B0(n90), .B1(sta25[1]), .C0(n108), 
        .C1(N405), .Y(n125) );
  OAI222XL U59 ( .A0(n63), .A1(n88), .B0(n72), .B1(n107), .C0(n97), .C1(n125), 
        .Y(N468) );
  AOI222XL U60 ( .A0(sta25[2]), .A1(n90), .B0(n99), .B1(sta21[2]), .C0(n108), 
        .C1(N406), .Y(n126) );
  OAI222XL U61 ( .A0(n62), .A1(n88), .B0(n71), .B1(n107), .C0(n97), .C1(n126), 
        .Y(N469) );
  OAI21XL U71 ( .A0(n133), .A1(n134), .B0(n135), .Y(n307) );
  OAI22XL U76 ( .A0(n146), .A1(n68), .B0(n69), .B1(n147), .Y(n145) );
  OAI22XL U77 ( .A0(n148), .A1(n68), .B0(n149), .B1(n80), .Y(n144) );
  OAI2BB1X1 U78 ( .A0N(sta26[1]), .A1N(n150), .B0(n151), .Y(n309) );
  OAI222XL U80 ( .A0(n66), .A1(n93), .B0(n147), .B1(sta26[1]), .C0(n81), .C1(
        n149), .Y(n152) );
  OAI21XL U82 ( .A0(n46), .A1(n146), .B0(n139), .Y(n150) );
  OAI222XL U84 ( .A0(n139), .A1(n70), .B0(n46), .B1(n156), .C0(n140), .C1(n157), .Y(n310) );
  OAI22XL U86 ( .A0(n154), .A1(n70), .B0(n82), .B1(n149), .Y(n158) );
  OAI22XL U96 ( .A0(n171), .A1(n65), .B0(n172), .B1(n68), .Y(n166) );
  OA22X1 U99 ( .A0(n175), .A1(n46), .B0(n66), .B1(n162), .Y(n173) );
  AOI222XL U100 ( .A0(n176), .A1(sta22[1]), .B0(n94), .B1(sta26[1]), .C0(n66), 
        .C1(n165), .Y(n175) );
  OAI222XL U102 ( .A0(n162), .A1(n67), .B0(n46), .B1(n177), .C0(n163), .C1(
        n157), .Y(n313) );
  OAI22XL U104 ( .A0(n92), .A1(n61), .B0(n70), .B1(n172), .Y(n178) );
  OAI31XL U106 ( .A0(n171), .A1(n66), .A2(n65), .B0(n179), .Y(n170) );
  OAI22XL U111 ( .A0(n187), .A1(n59), .B0(n60), .B1(n188), .Y(n186) );
  OAI22XL U113 ( .A0(n171), .A1(n59), .B0(n149), .B1(n65), .Y(n185) );
  OAI222XL U117 ( .A0(n66), .A1(n149), .B0(n188), .B1(sta22[1]), .C0(n81), 
        .C1(n93), .Y(n193) );
  OAI222XL U119 ( .A0(n182), .A1(n61), .B0(n46), .B1(n194), .C0(n183), .C1(
        n157), .Y(n316) );
  OAI22XL U121 ( .A0(n93), .A1(n82), .B0(n149), .B1(n67), .Y(n195) );
  OAI31XL U124 ( .A0(n171), .A1(n60), .A2(n59), .B0(n179), .Y(n190) );
  OA22X1 U130 ( .A0(n201), .A1(n86), .B0(n202), .B1(n142), .Y(n199) );
  AO22X1 U132 ( .A0(sta20[2]), .A1(n205), .B0(sta20[1]), .B1(n206), .Y(n204)
         );
  OAI22XL U133 ( .A0(n148), .A1(n80), .B0(n172), .B1(n59), .Y(n203) );
  OAI21XL U134 ( .A0(n201), .A1(n153), .B0(n207), .Y(n318) );
  OAI22XL U136 ( .A0(n209), .A1(n46), .B0(n81), .B1(n200), .Y(n208) );
  AOI222XL U137 ( .A0(n176), .A1(sta26[1]), .B0(n94), .B1(sta22[1]), .C0(n81), 
        .C1(n206), .Y(n209) );
  OAI222XL U140 ( .A0(n200), .A1(n82), .B0(n46), .B1(n212), .C0(n201), .C1(
        n157), .Y(n319) );
  OAI22XL U142 ( .A0(n211), .A1(n82), .B0(n172), .B1(n61), .Y(n213) );
  OAI2BB1X1 U145 ( .A0N(n95), .A1N(n197), .B0(n214), .Y(n159) );
  NAND3BX1 U147 ( .AN(mode[1]), .B(mode[0]), .C(mode[2]), .Y(n148) );
  OAI21XL U154 ( .A0(n216), .A1(n157), .B0(n217), .Y(n320) );
  OAI21XL U156 ( .A0(n216), .A1(n153), .B0(n219), .Y(n321) );
  OAI21XL U158 ( .A0(n216), .A1(n134), .B0(n220), .Y(n322) );
  NAND3BX1 U161 ( .AN(cnt1[1]), .B(cnt1[2]), .C(n221), .Y(n216) );
  OAI21XL U164 ( .A0(n47), .A1(n225), .B0(sta24[2]), .Y(n222) );
  OAI21XL U165 ( .A0(n54), .A1(n153), .B0(n227), .Y(n324) );
  OAI22XL U166 ( .A0(sta24[1]), .A1(n224), .B0(n75), .B1(n225), .Y(n227) );
  OAI21XL U167 ( .A0(sta24[0]), .A1(n226), .B0(n228), .Y(n225) );
  OAI222XL U169 ( .A0(n228), .A1(n76), .B0(n226), .B1(sta24[0]), .C0(n54), 
        .C1(n157), .Y(n325) );
  NAND3BX1 U177 ( .AN(mode[0]), .B(mode[2]), .C(mode[1]), .Y(n230) );
  OAI21XL U178 ( .A0(n233), .A1(n157), .B0(n234), .Y(n326) );
  OAI21XL U180 ( .A0(n233), .A1(n153), .B0(n236), .Y(n327) );
  OAI21XL U182 ( .A0(n233), .A1(n134), .B0(n237), .Y(n328) );
  OAI21XL U186 ( .A0(n238), .A1(n157), .B0(n239), .Y(n329) );
  OAI21XL U188 ( .A0(n238), .A1(n153), .B0(n241), .Y(n330) );
  OAI21XL U190 ( .A0(n238), .A1(n134), .B0(n242), .Y(n331) );
  AO22X1 U198 ( .A0(cnt1[17]), .A1(n244), .B0(n435), .B1(N70), .Y(n335) );
  AO22X1 U199 ( .A0(cnt1[16]), .A1(n244), .B0(n435), .B1(N69), .Y(n336) );
  AO22X1 U200 ( .A0(cnt1[15]), .A1(n244), .B0(n435), .B1(N68), .Y(n337) );
  AO22X1 U201 ( .A0(cnt1[14]), .A1(n244), .B0(n435), .B1(N67), .Y(n338) );
  AO22X1 U203 ( .A0(cnt1[12]), .A1(n244), .B0(n435), .B1(N65), .Y(n340) );
  AO22X1 U204 ( .A0(cnt1[11]), .A1(n244), .B0(n435), .B1(N64), .Y(n341) );
  AO22X1 U205 ( .A0(cnt1[10]), .A1(n244), .B0(n435), .B1(N63), .Y(n342) );
  AO22X1 U206 ( .A0(cnt1[9]), .A1(n244), .B0(n435), .B1(N62), .Y(n343) );
  AO22X1 U207 ( .A0(cnt1[8]), .A1(n244), .B0(n435), .B1(N61), .Y(n344) );
  AO22X1 U208 ( .A0(cnt1[7]), .A1(n244), .B0(n435), .B1(N60), .Y(n345) );
  AO22X1 U209 ( .A0(cnt1[6]), .A1(n244), .B0(n435), .B1(N59), .Y(n346) );
  AO22X1 U210 ( .A0(cnt1[5]), .A1(n244), .B0(n435), .B1(N58), .Y(n347) );
  AO22X1 U213 ( .A0(cnt1[2]), .A1(n244), .B0(n435), .B1(N55), .Y(n350) );
  AO22X1 U214 ( .A0(cnt1[1]), .A1(n244), .B0(n435), .B1(N54), .Y(n351) );
  AO22X1 U215 ( .A0(cnt1[0]), .A1(n244), .B0(n435), .B1(N53), .Y(n352) );
  AO22X1 U217 ( .A0(n44), .A1(n52), .B0(cnt2[0]), .B1(n245), .Y(n353) );
  AO22X1 U218 ( .A0(n44), .A1(N76), .B0(cnt2[1]), .B1(n245), .Y(n354) );
  AO22X1 U219 ( .A0(n44), .A1(N77), .B0(cnt2[2]), .B1(n245), .Y(n355) );
  AO22X1 U236 ( .A0(n44), .A1(N94), .B0(cnt2[19]), .B1(n245), .Y(n372) );
  OAI22XL U243 ( .A0(cnt2[3]), .A1(n252), .B0(n49), .B1(n50), .Y(n250) );
  OAI222XL U248 ( .A0(n76), .A1(n259), .B0(n79), .B1(n260), .C0(n61), .C1(n261), .Y(n258) );
  OAI22XL U250 ( .A0(n70), .A1(n265), .B0(n67), .B1(n266), .Y(n264) );
  OAI22XL U251 ( .A0(n82), .A1(n267), .B0(n85), .B1(n268), .Y(n263) );
  OAI22XL U255 ( .A0(n60), .A1(n261), .B0(n72), .B1(n257), .Y(n273) );
  OAI22XL U256 ( .A0(n75), .A1(n259), .B0(n78), .B1(n260), .Y(n272) );
  OAI22XL U258 ( .A0(n69), .A1(n265), .B0(n66), .B1(n266), .Y(n275) );
  OAI22XL U259 ( .A0(n81), .A1(n267), .B0(n84), .B1(n268), .Y(n274) );
  OAI31XL U260 ( .A0(n276), .A1(n253), .A2(n251), .B0(n277), .Y(n304) );
  OAI31XL U263 ( .A0(cnt2[1]), .A1(cnt2[2]), .A2(n49), .B0(n279), .Y(n278) );
  OAI31XL U264 ( .A0(cnt2[1]), .A1(cnt2[2]), .A2(cnt2[0]), .B0(n49), .Y(n279)
         );
  NOR3BXL U273 ( .AN(n285), .B(n286), .C(n287), .Y(n276) );
  OAI22XL U274 ( .A0(n59), .A1(n261), .B0(n71), .B1(n257), .Y(n287) );
  OAI22XL U277 ( .A0(n74), .A1(n259), .B0(n77), .B1(n260), .Y(n286) );
  OAI22XL U281 ( .A0(n68), .A1(n265), .B0(n65), .B1(n266), .Y(n291) );
  OAI22XL U284 ( .A0(n80), .A1(n267), .B0(n83), .B1(n268), .Y(n290) );
  OAI21XL U292 ( .A0(n133), .A1(n157), .B0(n293), .Y(n305) );
  OAI21XL U295 ( .A0(n133), .A1(n153), .B0(n294), .Y(n306) );
  NAND2BX1 U306 ( .AN(cnt1[3]), .B(n295), .Y(n180) );
  OAI21XL U314 ( .A0(n78), .A1(n79), .B0(n77), .Y(N450) );
  OAI2BB2XL U315 ( .B0(sta25[1]), .B1(N448), .A0N(sta25[1]), .A1N(N448), .Y(
        N449) );
  OAI21XL U316 ( .A0(n77), .A1(n78), .B0(sta25[0]), .Y(N448) );
  OAI21XL U317 ( .A0(n63), .A1(N433), .B0(n62), .Y(N435) );
  OAI2BB2XL U318 ( .B0(sta27[1]), .B1(N433), .A0N(sta27[1]), .A1N(N433), .Y(
        N434) );
  OAI21XL U319 ( .A0(n62), .A1(n63), .B0(sta27[0]), .Y(N433) );
  OAI21XL U320 ( .A0(n85), .A1(n84), .B0(n83), .Y(N421) );
  OAI2BB2XL U321 ( .B0(sta21[1]), .B1(N419), .A0N(sta21[1]), .A1N(N419), .Y(
        N420) );
  OAI21XL U322 ( .A0(n84), .A1(n83), .B0(sta21[0]), .Y(N419) );
  OAI21XL U323 ( .A0(n72), .A1(N404), .B0(n71), .Y(N406) );
  OAI2BB2XL U324 ( .B0(sta23[1]), .B1(N404), .A0N(sta23[1]), .A1N(N404), .Y(
        N405) );
  OAI21XL U325 ( .A0(n71), .A1(n72), .B0(sta23[0]), .Y(N404) );
  DFFRX1 sta10_reg_0_ ( .D(n319), .CK(clk), .RN(rst_n), .Q(sta20[0]), .QN(n82)
         );
  DFFRX1 sta15_reg_0_ ( .D(n320), .CK(clk), .RN(rst_n), .Q(sta25[0]), .QN(n79)
         );
  DFFRX1 sta14_reg_0_ ( .D(n325), .CK(clk), .RN(rst_n), .Q(sta24[0]), .QN(n76)
         );
  DFFRX1 sta_reg ( .D(n375), .CK(clk), .RN(rst_n), .Q(sta) );
  DFFRX1 sta13_reg_0_ ( .D(n326), .CK(clk), .RN(rst_n), .Q(sta23[0]), .QN(n73)
         );
  DFFRX1 sta12_reg_0_ ( .D(n316), .CK(clk), .RN(rst_n), .Q(sta22[0]), .QN(n61)
         );
  DFFRX1 sta16_reg_2_ ( .D(n308), .CK(clk), .RN(rst_n), .Q(sta26[2]), .QN(n68)
         );
  DFFRX1 sta11_reg_0_ ( .D(n305), .CK(clk), .RN(rst_n), .Q(sta21[0]), .QN(n85)
         );
  DFFRX1 cnt2_reg_20_ ( .D(n374), .CK(clk), .RN(rst_n), .Q(cnt2[20]) );
  DFFRX1 sta10_reg_1_ ( .D(n318), .CK(clk), .RN(rst_n), .Q(sta20[1]), .QN(n81)
         );
  DFFRX1 sta17_reg_2_ ( .D(n331), .CK(clk), .RN(rst_n), .Q(sta27[2]), .QN(n62)
         );
  DFFRX1 sta17_reg_1_ ( .D(n330), .CK(clk), .RN(rst_n), .Q(sta27[1]), .QN(n63)
         );
  DFFRX1 sta10_reg_2_ ( .D(n317), .CK(clk), .RN(rst_n), .Q(sta20[2]), .QN(n80)
         );
  DFFRX1 sta16_reg_0_ ( .D(n310), .CK(clk), .RN(rst_n), .Q(sta26[0]), .QN(n70)
         );
  DFFRX1 sta18_reg_0_ ( .D(n313), .CK(clk), .RN(rst_n), .Q(sta28[0]), .QN(n67)
         );
  DFFRX1 sta12_reg_1_ ( .D(n315), .CK(clk), .RN(rst_n), .Q(sta22[1]), .QN(n60)
         );
  DFFRX1 sta11_reg_2_ ( .D(n307), .CK(clk), .RN(rst_n), .Q(sta21[2]), .QN(n83)
         );
  DFFRX1 sta16_reg_1_ ( .D(n309), .CK(clk), .RN(rst_n), .Q(sta26[1]), .QN(n69)
         );
  DFFRX1 sta11_reg_1_ ( .D(n306), .CK(clk), .RN(rst_n), .Q(sta21[1]), .QN(n84)
         );
  DFFRX1 sta13_reg_2_ ( .D(n328), .CK(clk), .RN(rst_n), .Q(sta23[2]), .QN(n71)
         );
  DFFRX1 sta13_reg_1_ ( .D(n327), .CK(clk), .RN(rst_n), .Q(sta23[1]), .QN(n72)
         );
  DFFRX1 sta18_reg_2_ ( .D(n311), .CK(clk), .RN(rst_n), .Q(sta28[2]), .QN(n65)
         );
  DFFRX1 sta18_reg_1_ ( .D(n312), .CK(clk), .RN(rst_n), .Q(sta28[1]), .QN(n66)
         );
  DFFRX1 sta12_reg_2_ ( .D(n314), .CK(clk), .RN(rst_n), .QN(n59) );
  DFFRX1 sta17_reg_0_ ( .D(n329), .CK(clk), .RN(rst_n), .Q(sta27[0]), .QN(n64)
         );
  DFFRX1 sta14_reg_2_ ( .D(n323), .CK(clk), .RN(rst_n), .Q(sta24[2]), .QN(n74)
         );
  DFFRX1 sta15_reg_2_ ( .D(n322), .CK(clk), .RN(rst_n), .Q(sta25[2]), .QN(n77)
         );
  DFFRX1 sta15_reg_1_ ( .D(n321), .CK(clk), .RN(rst_n), .Q(sta25[1]), .QN(n78)
         );
  DFFRX1 sta14_reg_1_ ( .D(n324), .CK(clk), .RN(rst_n), .Q(sta24[1]), .QN(n75)
         );
  DFFRX1 cnt2_reg_18_ ( .D(n371), .CK(clk), .RN(rst_n), .Q(cnt2[18]) );
  DFFRX1 cnt2_reg_13_ ( .D(n366), .CK(clk), .RN(rst_n), .Q(cnt2[13]) );
  DFFRX1 cnt2_reg_17_ ( .D(n370), .CK(clk), .RN(rst_n), .Q(cnt2[17]) );
  DFFRX1 cnt2_reg_15_ ( .D(n368), .CK(clk), .RN(rst_n), .Q(cnt2[15]) );
  DFFRX1 cnt2_reg_16_ ( .D(n369), .CK(clk), .RN(rst_n), .Q(cnt2[16]) );
  DFFRX1 cnt2_reg_14_ ( .D(n367), .CK(clk), .RN(rst_n), .Q(cnt2[14]) );
  DFFRX1 cnt2_reg_9_ ( .D(n362), .CK(clk), .RN(rst_n), .Q(cnt2[9]) );
  DFFRX1 cnt1_reg_12_ ( .D(n340), .CK(clk), .RN(rst_n), .Q(cnt1[12]) );
  DFFRX1 cnt2_reg_7_ ( .D(n360), .CK(clk), .RN(rst_n), .Q(cnt2[7]) );
  DFFRX1 cnt2_reg_11_ ( .D(n364), .CK(clk), .RN(rst_n), .Q(cnt2[11]) );
  DFFRX1 cnt2_reg_8_ ( .D(n361), .CK(clk), .RN(rst_n), .Q(cnt2[8]) );
  DFFRX1 cnt2_reg_12_ ( .D(n365), .CK(clk), .RN(rst_n), .Q(cnt2[12]) );
  DFFRX1 cnt2_reg_6_ ( .D(n359), .CK(clk), .RN(rst_n), .Q(cnt2[6]) );
  DFFRX1 cnt2_reg_10_ ( .D(n363), .CK(clk), .RN(rst_n), .Q(cnt2[10]) );
  DFFRX1 out_valid_reg ( .D(n301), .CK(clk), .RN(rst_n), .Q(out_valid) );
  DFFRX1 out_reg_1_ ( .D(n303), .CK(clk), .RN(rst_n), .Q(out[1]) );
  DFFRX1 out_reg_0_ ( .D(n302), .CK(clk), .RN(rst_n), .Q(out[0]) );
  DFFRX1 out_reg_2_ ( .D(n304), .CK(clk), .RN(rst_n), .Q(out[2]) );
  DFFRX1 rst_reg ( .D(n373), .CK(clk), .RN(rst_n), .Q(rst), .QN(n45) );
  DFFRX1 cnt1_reg_20_ ( .D(n332), .CK(clk), .RN(rst_n), .Q(cnt1[20]) );
  DFFRX1 cnt2_reg_5_ ( .D(n358), .CK(clk), .RN(rst_n), .Q(cnt2[5]) );
  DFFRX1 cnt2_reg_4_ ( .D(n357), .CK(clk), .RN(rst_n), .Q(cnt2[4]) );
  DFFRX1 cnt1_reg_10_ ( .D(n342), .CK(clk), .RN(rst_n), .Q(cnt1[10]) );
  DFFRX1 cnt1_reg_11_ ( .D(n341), .CK(clk), .RN(rst_n), .Q(cnt1[11]) );
  DFFRX1 cnt1_reg_9_ ( .D(n343), .CK(clk), .RN(rst_n), .Q(cnt1[9]) );
  DFFRX1 cnt1_reg_7_ ( .D(n345), .CK(clk), .RN(rst_n), .Q(cnt1[7]) );
  DFFRX1 cnt1_reg_17_ ( .D(n335), .CK(clk), .RN(rst_n), .Q(cnt1[17]) );
  DFFRX1 cnt1_reg_4_ ( .D(n348), .CK(clk), .RN(rst_n), .Q(cnt1[4]) );
  DFFRX1 cnt1_reg_15_ ( .D(n337), .CK(clk), .RN(rst_n), .Q(cnt1[15]) );
  DFFRX1 cnt1_reg_6_ ( .D(n346), .CK(clk), .RN(rst_n), .Q(cnt1[6]) );
  DFFRX1 cnt1_reg_18_ ( .D(n334), .CK(clk), .RN(rst_n), .Q(cnt1[18]) );
  DFFRX1 cnt1_reg_14_ ( .D(n338), .CK(clk), .RN(rst_n), .Q(cnt1[14]) );
  DFFRX1 cnt1_reg_5_ ( .D(n347), .CK(clk), .RN(rst_n), .Q(cnt1[5]) );
  DFFRX1 cnt1_reg_16_ ( .D(n336), .CK(clk), .RN(rst_n), .Q(cnt1[16]) );
  DFFRX1 cnt1_reg_8_ ( .D(n344), .CK(clk), .RN(rst_n), .Q(cnt1[8]) );
  DFFRX1 cnt1_reg_3_ ( .D(n349), .CK(clk), .RN(rst_n), .Q(cnt1[3]) );
  DFFRX1 cnt1_reg_2_ ( .D(n350), .CK(clk), .RN(rst_n), .Q(cnt1[2]), .QN(n57)
         );
  AOI32XL U107 ( .A0(n56), .A1(n45), .A2(n163), .B0(n98), .B1(n45), .Y(n162)
         );
  NAND3XL U128 ( .A(cnt1[1]), .B(n160), .C(n57), .Y(n183) );
  AOI32XL U127 ( .A0(n183), .A1(n45), .A2(n142), .B0(n98), .B1(n45), .Y(n182)
         );
  AOI211XL U171 ( .A0(n229), .A1(in_valid), .B0(rst), .C0(n136), .Y(n232) );
  NAND3XL U90 ( .A(cnt1[2]), .B(cnt1[1]), .C(n160), .Y(n140) );
  AOI32XL U89 ( .A0(n140), .A1(n45), .A2(n142), .B0(n98), .B1(n45), .Y(n139)
         );
  AOI32XL U152 ( .A0(n201), .A1(n45), .A2(n142), .B0(n98), .B1(n45), .Y(n200)
         );
  OAI211XL U160 ( .A0(n216), .A1(n98), .B0(n45), .C0(n46), .Y(n218) );
  NAND3XL U194 ( .A(cnt1[2]), .B(cnt1[1]), .C(n221), .Y(n238) );
  AOI211XL U192 ( .A0(n53), .A1(in_valid), .B0(rst), .C0(n136), .Y(n240) );
  AOI22XL U187 ( .A0(n136), .A1(N479), .B0(n240), .B1(sta27[0]), .Y(n239) );
  AOI22XL U189 ( .A0(n136), .A1(N480), .B0(n240), .B1(sta27[1]), .Y(n241) );
  AOI22XL U191 ( .A0(n136), .A1(N481), .B0(n240), .B1(sta27[2]), .Y(n242) );
  OAI211XL U184 ( .A0(n233), .A1(n98), .B0(n45), .C0(n46), .Y(n235) );
  OAI211XL U297 ( .A0(n133), .A1(n98), .B0(n45), .C0(n46), .Y(n137) );
  NAND3XL U283 ( .A(cnt2[1]), .B(cnt2[2]), .C(n289), .Y(n265) );
  NAND3XL U282 ( .A(cnt2[0]), .B(cnt2[3]), .C(n292), .Y(n266) );
  NAND3XL U278 ( .A(cnt2[1]), .B(cnt2[2]), .C(n288), .Y(n260) );
  AOI211XL U253 ( .A0(n270), .A1(n271), .B0(n253), .C0(n251), .Y(n269) );
  AOI211XL U246 ( .A0(n255), .A1(n256), .B0(n253), .C0(n251), .Y(n254) );
  NAND2XL U261 ( .A(n253), .B(out[2]), .Y(n277) );
  NAND4XL U238 ( .A(cnt2[3]), .B(n248), .C(n45), .D(n52), .Y(n247) );
  NOR2X1 U301 ( .A(cnt1[0]), .B(n180), .Y(n160) );
  NAND3X1 U308 ( .A(n298), .B(n299), .C(n300), .Y(n297) );
  CLKINVX1 U12 ( .A(in[2]), .Y(n86) );
  NAND3X1 U126 ( .A(mode[2]), .B(mode[1]), .C(mode[0]), .Y(n171) );
  NOR2X1 U101 ( .A(n171), .B(n67), .Y(n165) );
  NAND2X1 U143 ( .A(mode[0]), .B(n95), .Y(n172) );
  NAND2X1 U151 ( .A(mode[1]), .B(n95), .Y(n149) );
  NOR2X1 U150 ( .A(mode[1]), .B(mode[0]), .Y(n197) );
  NAND2X1 U149 ( .A(mode[2]), .B(n197), .Y(n196) );
  NOR2X1 U105 ( .A(sta28[0]), .B(n171), .Y(n169) );
  NAND2X1 U176 ( .A(mode[2]), .B(mode[1]), .Y(n214) );
  NOR2X1 U175 ( .A(mode[0]), .B(n214), .Y(n198) );
  AOI211X1 U125 ( .A0(n197), .A1(n95), .B0(n91), .C0(n198), .Y(n179) );
  AOI211X1 U93 ( .A0(sta28[1]), .A1(n165), .B0(n166), .C0(n167), .Y(n164) );
  NOR2X1 U123 ( .A(sta22[0]), .B(n171), .Y(n189) );
  AOI211X1 U110 ( .A0(sta20[2]), .A1(n143), .B0(n185), .C0(n186), .Y(n184) );
  NOR2X1 U168 ( .A(n76), .B(n226), .Y(n224) );
  AOI211X1 U170 ( .A0(n230), .A1(n136), .B0(n231), .C0(n232), .Y(n228) );
  NAND2X1 U163 ( .A(sta24[1]), .B(n224), .Y(n223) );
  AOI31X1 U87 ( .A0(n91), .A1(sta26[1]), .A2(sta26[2]), .B0(n159), .Y(n154) );
  NOR2X1 U88 ( .A(sta26[0]), .B(n148), .Y(n155) );
  NOR2BX1 U83 ( .AN(n154), .B(n155), .Y(n146) );
  AOI211X1 U75 ( .A0(sta28[2]), .A1(n143), .B0(n144), .C0(n145), .Y(n141) );
  NOR2X1 U146 ( .A(sta20[0]), .B(n148), .Y(n210) );
  AOI31X1 U144 ( .A0(n91), .A1(sta20[2]), .A2(sta20[1]), .B0(n159), .Y(n211)
         );
  NAND2BX1 U139 ( .AN(n210), .B(n211), .Y(n205) );
  AOI211X1 U131 ( .A0(sta26[2]), .A1(n176), .B0(n203), .C0(n204), .Y(n202) );
  NOR2X1 U34 ( .A(mode[1]), .B(n95), .Y(n108) );
  NAND2X1 U27 ( .A(mode[2]), .B(n97), .Y(n101) );
  NOR2X1 U30 ( .A(mode[1]), .B(n101), .Y(n104) );
  CLKINVX1 U22 ( .A(mode[1]), .Y(n96) );
  NOR2X1 U37 ( .A(n95), .B(n96), .Y(n111) );
  CLKINVX1 U15 ( .A(n109), .Y(n89) );
  CLKINVX1 U14 ( .A(n104), .Y(n88) );
  NOR2X1 U28 ( .A(n96), .B(n101), .Y(n102) );
  NAND2X1 U26 ( .A(mode[0]), .B(n99), .Y(n100) );
  AOI22X1 U65 ( .A0(n102), .A1(N420), .B0(n103), .B1(sta27[1]), .Y(n129) );
  AOI22X1 U62 ( .A0(n102), .A1(N419), .B0(n103), .B1(sta27[0]), .Y(n127) );
  AOI22X1 U68 ( .A0(n102), .A1(N421), .B0(sta27[2]), .B1(n103), .Y(n131) );
  OAI211X1 U70 ( .A0(n77), .A1(n100), .B0(n131), .C0(n132), .Y(N463) );
  NAND4X1 U266 ( .A(n280), .B(n281), .C(n282), .D(n283), .Y(n246) );
  NOR2X1 U289 ( .A(cnt2[3]), .B(n52), .Y(n289) );
  AOI211X1 U257 ( .A0(sta27[1]), .A1(n262), .B0(n274), .C0(n275), .Y(n270) );
  AOI211X1 U249 ( .A0(sta27[0]), .A1(n262), .B0(n263), .C0(n264), .Y(n255) );
  NAND2X1 U193 ( .A(n435), .B(in[2]), .Y(n134) );
  OAI22XL U73 ( .A0(n138), .A1(n434), .B0(n68), .B1(n139), .Y(n308) );
  NAND3XL U185 ( .A(cnt1[1]), .B(n221), .C(n57), .Y(n233) );
  AOI31XL U135 ( .A0(n136), .A1(sta20[1]), .A2(n205), .B0(n208), .Y(n207) );
  NAND3XL U279 ( .A(cnt2[2]), .B(n289), .C(n51), .Y(n259) );
  OAI22XL U108 ( .A0(n181), .A1(n434), .B0(n59), .B1(n182), .Y(n314) );
  NOR3XL U172 ( .A(n57), .B(n55), .C(cnt1[1]), .Y(n229) );
  OAI22XL U129 ( .A0(n199), .A1(n434), .B0(n80), .B1(n200), .Y(n317) );
  OAI211XL U98 ( .A0(n169), .A1(n170), .B0(sta28[1]), .C0(n136), .Y(n174) );
  OAI211XL U115 ( .A0(n189), .A1(n190), .B0(sta22[1]), .C0(n136), .Y(n192) );
  NOR4XL U271 ( .A(cnt2[6]), .B(cnt2[7]), .C(cnt2[8]), .D(cnt2[9]), .Y(n280)
         );
  NOR4XL U270 ( .A(cnt2[10]), .B(cnt2[11]), .C(cnt2[12]), .D(cnt2[13]), .Y(
        n281) );
  NOR4XL U269 ( .A(cnt2[14]), .B(cnt2[15]), .C(cnt2[16]), .D(cnt2[17]), .Y(
        n282) );
  NAND3XL U275 ( .A(cnt2[2]), .B(n288), .C(n51), .Y(n257) );
  NOR2XL U313 ( .A(cnt1[2]), .B(cnt1[1]), .Y(n215) );
  NOR2XL U291 ( .A(cnt2[1]), .B(cnt2[2]), .Y(n292) );
  NOR2XL U287 ( .A(cnt2[0]), .B(cnt2[3]), .Y(n288) );
  NOR3X1 U307 ( .A(cnt1[12]), .B(n296), .C(n297), .Y(n295) );
  NOR2XL U286 ( .A(cnt2[2]), .B(n51), .Y(n248) );
  AOI211XL U103 ( .A0(sta28[0]), .A1(n170), .B0(n169), .C0(n178), .Y(n177) );
  OR4X1 U312 ( .A(cnt1[11]), .B(cnt1[10]), .C(cnt1[7]), .D(cnt1[9]), .Y(n296)
         );
  AOI211XL U120 ( .A0(sta22[0]), .A1(n190), .B0(n189), .C0(n195), .Y(n194) );
  NOR2XL U138 ( .A(n148), .B(n82), .Y(n206) );
  OAI22XL U94 ( .A0(n92), .A1(n59), .B0(n168), .B1(n65), .Y(n167) );
  OAI22XL U91 ( .A0(n161), .A1(n434), .B0(n65), .B1(n162), .Y(n311) );
  DFFRX4 cnt2_reg_0_ ( .D(n353), .CK(clk), .RN(rst_n), .Q(cnt2[0]), .QN(n52)
         );
  DFFRX4 cnt2_reg_1_ ( .D(n354), .CK(clk), .RN(rst_n), .Q(cnt2[1]), .QN(n51)
         );
  DFFRX2 cnt2_reg_2_ ( .D(n355), .CK(clk), .RN(rst_n), .Q(cnt2[2]) );
  DFFRX2 cnt2_reg_3_ ( .D(n356), .CK(clk), .RN(rst_n), .Q(cnt2[3]), .QN(n49)
         );
  ADDHXL add_x_41_1_U1_1_18 ( .A(cnt2[18]), .B(add_x_41_1_carry_18_), .CO(
        add_x_41_1_carry_19_), .S(N93) );
  ADDHXL add_x_41_1_U1_1_17 ( .A(cnt2[17]), .B(add_x_41_1_carry_17_), .CO(
        add_x_41_1_carry_18_), .S(N92) );
  ADDHXL add_x_41_1_U1_1_16 ( .A(cnt2[16]), .B(add_x_41_1_carry_16_), .CO(
        add_x_41_1_carry_17_), .S(N91) );
  ADDHXL add_x_41_1_U1_1_11 ( .A(cnt2[11]), .B(add_x_41_1_carry_11_), .CO(
        add_x_41_1_carry_12_), .S(N86) );
  ADDHXL add_x_41_1_U1_1_10 ( .A(cnt2[10]), .B(add_x_41_1_carry_10_), .CO(
        add_x_41_1_carry_11_), .S(N85) );
  ADDHXL add_x_41_1_U1_1_9 ( .A(cnt2[9]), .B(add_x_41_1_carry_9_), .CO(
        add_x_41_1_carry_10_), .S(N84) );
  ADDHXL add_x_41_1_U1_1_8 ( .A(cnt2[8]), .B(add_x_41_1_carry_8_), .CO(
        add_x_41_1_carry_9_), .S(N83) );
  ADDHXL add_x_41_1_U1_1_7 ( .A(cnt2[7]), .B(add_x_41_1_carry_7_), .CO(
        add_x_41_1_carry_8_), .S(N82) );
  ADDHXL add_x_41_1_U1_1_6 ( .A(cnt2[6]), .B(add_x_41_1_carry_6_), .CO(
        add_x_41_1_carry_7_), .S(N81) );
  ADDHXL add_x_41_1_U1_1_5 ( .A(cnt2[5]), .B(add_x_41_1_carry_5_), .CO(
        add_x_41_1_carry_6_), .S(N80) );
  ADDHXL add_x_41_1_U1_1_4 ( .A(cnt2[4]), .B(add_x_41_1_carry_4_), .CO(
        add_x_41_1_carry_5_), .S(N79) );
  ADDHXL add_x_41_0_U1_1_17 ( .A(cnt1[17]), .B(add_x_41_0_carry_17_), .CO(
        add_x_41_0_carry_18_), .S(N70) );
  ADDHXL add_x_41_0_U1_1_16 ( .A(cnt1[16]), .B(add_x_41_0_carry_16_), .CO(
        add_x_41_0_carry_17_), .S(N69) );
  ADDHXL add_x_41_0_U1_1_15 ( .A(cnt1[15]), .B(add_x_41_0_carry_15_), .CO(
        add_x_41_0_carry_16_), .S(N68) );
  ADDHXL add_x_41_0_U1_1_12 ( .A(cnt1[12]), .B(add_x_41_0_carry_12_), .CO(
        add_x_41_0_carry_13_), .S(N65) );
  ADDHXL add_x_41_0_U1_1_11 ( .A(cnt1[11]), .B(add_x_41_0_carry_11_), .CO(
        add_x_41_0_carry_12_), .S(N64) );
  ADDHXL add_x_41_0_U1_1_10 ( .A(cnt1[10]), .B(add_x_41_0_carry_10_), .CO(
        add_x_41_0_carry_11_), .S(N63) );
  ADDHXL add_x_41_0_U1_1_9 ( .A(cnt1[9]), .B(add_x_41_0_carry_9_), .CO(
        add_x_41_0_carry_10_), .S(N62) );
  ADDHXL add_x_41_0_U1_1_8 ( .A(cnt1[8]), .B(add_x_41_0_carry_8_), .CO(
        add_x_41_0_carry_9_), .S(N61) );
  ADDHXL add_x_41_0_U1_1_7 ( .A(cnt1[7]), .B(add_x_41_0_carry_7_), .CO(
        add_x_41_0_carry_8_), .S(N60) );
  ADDHXL add_x_41_0_U1_1_6 ( .A(cnt1[6]), .B(add_x_41_0_carry_6_), .CO(
        add_x_41_0_carry_7_), .S(N59) );
  NAND2XL U31 ( .A(n95), .B(n96), .Y(n105) );
  NOR4X1 U310 ( .A(cnt1[20]), .B(cnt1[19]), .C(cnt1[18]), .D(cnt1[17]), .Y(
        n299) );
  NOR4X1 U311 ( .A(cnt1[8]), .B(cnt1[6]), .C(cnt1[5]), .D(cnt1[4]), .Y(n298)
         );
  NOR4X1 U309 ( .A(cnt1[16]), .B(cnt1[15]), .C(cnt1[14]), .D(cnt1[13]), .Y(
        n300) );
  OR2XL U118 ( .A(n171), .B(n61), .Y(n188) );
  OR4XL U268 ( .A(cnt2[19]), .B(cnt2[20]), .C(cnt2[4]), .D(cnt2[5]), .Y(n284)
         );
  INVXL U20 ( .A(n172), .Y(n94) );
  INVX1 U16 ( .A(n105), .Y(n90) );
  NAND2XL U81 ( .A(n91), .B(sta26[0]), .Y(n147) );
  NAND2XL U276 ( .A(n289), .B(n248), .Y(n261) );
  INVX1 U7 ( .A(n292), .Y(n50) );
  NOR2XL U267 ( .A(cnt2[18]), .B(n284), .Y(n283) );
  NAND2XL U285 ( .A(n288), .B(n248), .Y(n268) );
  NAND2XL U288 ( .A(n289), .B(n292), .Y(n267) );
  OAI2BB1XL U240 ( .A0N(sta), .A1N(n45), .B0(n434), .Y(n375) );
  AOI22XL U41 ( .A0(n99), .A1(n113), .B0(sta27[0]), .B1(n114), .Y(n115) );
  AOI22XL U47 ( .A0(n99), .A1(n110), .B0(sta27[2]), .B1(n114), .Y(n119) );
  AOI22XL U44 ( .A0(n99), .A1(n112), .B0(sta27[1]), .B1(n114), .Y(n117) );
  AOI22XL U69 ( .A0(n104), .A1(sta23[2]), .B0(sta21[2]), .B1(n106), .Y(n132)
         );
  AOI22XL U63 ( .A0(n104), .A1(sta23[0]), .B0(sta21[0]), .B1(n106), .Y(n128)
         );
  AOI22XL U66 ( .A0(n104), .A1(sta23[1]), .B0(sta21[1]), .B1(n106), .Y(n130)
         );
  NAND2XL U42 ( .A(n102), .B(N433), .Y(n116) );
  NOR2XL U244 ( .A(cnt2[0]), .B(n50), .Y(n252) );
  NAND2XL U48 ( .A(n102), .B(N435), .Y(n120) );
  NAND2XL U45 ( .A(n102), .B(N434), .Y(n118) );
  NOR3X1 U290 ( .A(cnt2[0]), .B(n49), .C(n50), .Y(n262) );
  NOR2XL U112 ( .A(n189), .B(n190), .Y(n187) );
  AOI211XL U141 ( .A0(sta26[0]), .A1(n176), .B0(n210), .C0(n213), .Y(n212) );
  AOI211XL U85 ( .A0(sta28[0]), .A1(n143), .B0(n155), .C0(n158), .Y(n156) );
  NOR2XL U95 ( .A(n169), .B(n170), .Y(n168) );
  OAI211XL U43 ( .A0(n79), .A1(n88), .B0(n115), .C0(n116), .Y(N479) );
  NOR2XL U237 ( .A(n246), .B(n247), .Y(n373) );
  NOR2XL U265 ( .A(n251), .B(n246), .Y(n249) );
  NAND4X1 U300 ( .A(n215), .B(cnt1[3]), .C(n295), .D(N53), .Y(n163) );
  NOR2XL U254 ( .A(n272), .B(n273), .Y(n271) );
  AOI211XL U280 ( .A0(sta27[2]), .A1(n262), .B0(n290), .C0(n291), .Y(n285) );
  AO22XL U220 ( .A0(n44), .A1(N78), .B0(cnt2[3]), .B1(n245), .Y(n356) );
  OAI211XL U49 ( .A0(n88), .A1(n77), .B0(n119), .C0(n120), .Y(N481) );
  AOI2BB1XL U247 ( .A0N(n257), .A1N(n73), .B0(n258), .Y(n256) );
  OAI211XL U46 ( .A0(n78), .A1(n88), .B0(n117), .C0(n118), .Y(N480) );
  OAI211XL U67 ( .A0(n100), .A1(n78), .B0(n129), .C0(n130), .Y(N462) );
  OAI211XL U64 ( .A0(n100), .A1(n79), .B0(n127), .C0(n128), .Y(N461) );
  AO22XL U221 ( .A0(n44), .A1(N79), .B0(cnt2[4]), .B1(n245), .Y(n357) );
  NOR2X1 U305 ( .A(N53), .B(n180), .Y(n221) );
  AO22XL U241 ( .A0(n249), .A1(n250), .B0(n245), .B1(out_valid), .Y(n301) );
  INVXL U11 ( .A(n180), .Y(n56) );
  AOI21X1 U262 ( .A0(n249), .A1(n278), .B0(rst), .Y(n253) );
  AO22XL U222 ( .A0(n44), .A1(N80), .B0(cnt2[5]), .B1(n245), .Y(n358) );
  NAND2XL U153 ( .A(n215), .B(n160), .Y(n201) );
  NAND2XL U304 ( .A(n215), .B(n221), .Y(n133) );
  INVX1 U10 ( .A(n160), .Y(n55) );
  AO21XL U245 ( .A0(n253), .A1(out[0]), .B0(n254), .Y(n302) );
  AO22XL U223 ( .A0(n44), .A1(N81), .B0(cnt2[6]), .B1(n245), .Y(n359) );
  AO21XL U252 ( .A0(n253), .A1(out[1]), .B0(n269), .Y(n303) );
  INVXL U8 ( .A(n238), .Y(n53) );
  OA22XL U74 ( .A0(n140), .A1(n86), .B0(n141), .B1(n142), .Y(n138) );
  OA22XL U109 ( .A0(n183), .A1(n86), .B0(n184), .B1(n142), .Y(n181) );
  INVX1 U9 ( .A(n229), .Y(n54) );
  OA22XL U92 ( .A0(n163), .A1(n86), .B0(n164), .B1(n142), .Y(n161) );
  AO22XL U224 ( .A0(n44), .A1(N82), .B0(cnt2[7]), .B1(n245), .Y(n360) );
  AO22XL U225 ( .A0(n44), .A1(N83), .B0(cnt2[8]), .B1(n245), .Y(n361) );
  AOI2BB2XL U116 ( .B0(n136), .B1(n193), .A0N(n60), .A1N(n182), .Y(n191) );
  AOI2BB2XL U79 ( .B0(n136), .B1(n152), .A0N(n153), .A1N(n140), .Y(n151) );
  OAI211XL U114 ( .A0(n153), .A1(n183), .B0(n191), .C0(n192), .Y(n315) );
  AO22XL U226 ( .A0(n44), .A1(N84), .B0(cnt2[9]), .B1(n245), .Y(n362) );
  INVXL U5 ( .A(n226), .Y(n47) );
  AOI2BB2XL U183 ( .B0(n136), .B1(N469), .A0N(n235), .A1N(n71), .Y(n237) );
  AOI2BB2XL U157 ( .B0(n136), .B1(N474), .A0N(n218), .A1N(n78), .Y(n219) );
  OAI211XL U97 ( .A0(n153), .A1(n163), .B0(n173), .C0(n174), .Y(n312) );
  AOI2BB2XL U181 ( .B0(n136), .B1(N468), .A0N(n235), .A1N(n72), .Y(n236) );
  AOI2BB2XL U72 ( .B0(n136), .B1(N463), .A0N(n137), .A1N(n83), .Y(n135) );
  AOI2BB2XL U159 ( .B0(n136), .B1(N475), .A0N(n218), .A1N(n77), .Y(n220) );
  AOI2BB2XL U293 ( .B0(n136), .B1(N461), .A0N(n137), .A1N(n85), .Y(n293) );
  AO22XL U227 ( .A0(n44), .A1(N85), .B0(cnt2[10]), .B1(n245), .Y(n363) );
  AOI2BB2XL U296 ( .B0(n136), .B1(N462), .A0N(n137), .A1N(n84), .Y(n294) );
  AOI2BB2XL U155 ( .B0(n136), .B1(N473), .A0N(n218), .A1N(n79), .Y(n217) );
  AOI2BB2XL U179 ( .B0(n136), .B1(N467), .A0N(n235), .A1N(n73), .Y(n234) );
  AO22XL U228 ( .A0(n44), .A1(N86), .B0(cnt2[11]), .B1(n245), .Y(n364) );
  AO22XL U229 ( .A0(n44), .A1(N87), .B0(cnt2[12]), .B1(n245), .Y(n365) );
  OAI211XL U162 ( .A0(n134), .A1(n54), .B0(n222), .C0(n223), .Y(n323) );
  AO22XL U230 ( .A0(n44), .A1(N88), .B0(cnt2[13]), .B1(n245), .Y(n366) );
  AO22XL U231 ( .A0(n44), .A1(N89), .B0(cnt2[14]), .B1(n245), .Y(n367) );
  AO22XL U232 ( .A0(n44), .A1(N90), .B0(cnt2[15]), .B1(n245), .Y(n368) );
  AO22XL U233 ( .A0(n44), .A1(N91), .B0(cnt2[16]), .B1(n245), .Y(n369) );
  AO22XL U234 ( .A0(n44), .A1(N92), .B0(cnt2[17]), .B1(n245), .Y(n370) );
  AO22XL U235 ( .A0(n44), .A1(N93), .B0(cnt2[18]), .B1(n245), .Y(n371) );
  DFFRHQX2 cnt1_reg_1_ ( .D(n351), .CK(clk), .RN(rst_n), .Q(cnt1[1]) );
  DFFRX1 cnt1_reg_0_ ( .D(n352), .CK(clk), .RN(rst_n), .Q(cnt1[0]), .QN(N53)
         );
  DFFRX1 cnt1_reg_19_ ( .D(n333), .CK(clk), .RN(rst_n), .Q(cnt1[19]) );
  DFFRX2 cnt2_reg_19_ ( .D(n372), .CK(clk), .RN(rst_n), .Q(cnt2[19]) );
  DFFRX1 cnt1_reg_13_ ( .D(n339), .CK(clk), .RN(rst_n), .Q(cnt1[13]) );
  CLKINVX1 U327 ( .A(1'b0), .Y(ready) );
  CLKINVX1 U329 ( .A(mode[2]), .Y(n95) );
  INVX3 U330 ( .A(in_valid), .Y(n98) );
  ADDHXL U331 ( .A(cnt1[1]), .B(cnt1[0]), .CO(add_x_41_0_carry_2_), .S(N54) );
  AND2X2 U332 ( .A(cnt1[3]), .B(add_x_41_0_carry_3_), .Y(n391) );
  AND2X2 U333 ( .A(cnt1[18]), .B(add_x_41_0_carry_18_), .Y(n392) );
  NAND3X1 U334 ( .A(sta), .B(n45), .C(n98), .Y(n251) );
  CLKINVX1 U335 ( .A(n434), .Y(n435) );
  NOR2X1 U336 ( .A(rst), .B(in_valid), .Y(n244) );
  NAND2X1 U337 ( .A(n435), .B(in[1]), .Y(n153) );
  NAND2X1 U338 ( .A(cnt2[19]), .B(add_x_41_1_carry_19_), .Y(n394) );
  NOR2X1 U339 ( .A(rst), .B(n44), .Y(n245) );
  CLKINVX1 U340 ( .A(n251), .Y(n44) );
  OAI21XL U341 ( .A0(mode[1]), .A1(n172), .B0(n196), .Y(n143) );
  NAND3BX1 U342 ( .AN(n221), .B(n55), .C(n163), .Y(n142) );
  NOR2X1 U343 ( .A(n142), .B(n434), .Y(n136) );
  OAI21XL U344 ( .A0(mode[0]), .A1(n149), .B0(n196), .Y(n176) );
  CLKINVX1 U345 ( .A(n136), .Y(n46) );
  NAND2X1 U346 ( .A(n435), .B(in[0]), .Y(n157) );
  NOR3BX1 U347 ( .AN(cnt1[1]), .B(n57), .C(N53), .Y(add_x_41_0_carry_3_) );
  AOI2BB2X1 U348 ( .B0(cnt1[13]), .B1(add_x_41_0_carry_13_), .A0N(cnt1[13]), 
        .A1N(add_x_41_0_carry_13_), .Y(n381) );
  AO22X1 U349 ( .A0(cnt1[13]), .A1(n244), .B0(n381), .B1(n435), .Y(n339) );
  AND3X1 U350 ( .A(n391), .B(cnt1[4]), .C(cnt1[5]), .Y(add_x_41_0_carry_6_) );
  AND2X1 U351 ( .A(n391), .B(cnt1[4]), .Y(n382) );
  AOI2BB2X1 U352 ( .B0(n382), .B1(cnt1[5]), .A0N(n382), .A1N(cnt1[5]), .Y(N58)
         );
  AOI2BB2X1 U353 ( .B0(cnt1[19]), .B1(n392), .A0N(cnt1[19]), .A1N(n392), .Y(
        n383) );
  AO22X1 U354 ( .A0(cnt1[19]), .A1(n244), .B0(n383), .B1(n435), .Y(n333) );
  XOR2X1 U355 ( .A(cnt1[2]), .B(add_x_41_0_carry_2_), .Y(N55) );
  AOI2BB2X1 U356 ( .B0(cnt1[18]), .B1(add_x_41_0_carry_18_), .A0N(cnt1[18]), 
        .A1N(add_x_41_0_carry_18_), .Y(n384) );
  AO22X1 U357 ( .A0(cnt1[18]), .A1(n244), .B0(n384), .B1(n435), .Y(n334) );
  AOI2BB2X1 U358 ( .B0(cnt1[4]), .B1(n391), .A0N(cnt1[4]), .A1N(n391), .Y(n385) );
  AO22X1 U359 ( .A0(cnt1[4]), .A1(n244), .B0(n385), .B1(n435), .Y(n348) );
  AND3X1 U360 ( .A(add_x_41_0_carry_13_), .B(cnt1[13]), .C(cnt1[14]), .Y(
        add_x_41_0_carry_15_) );
  AND2X1 U361 ( .A(add_x_41_0_carry_13_), .B(cnt1[13]), .Y(n386) );
  AOI2BB2X1 U362 ( .B0(n386), .B1(cnt1[14]), .A0N(n386), .A1N(cnt1[14]), .Y(
        N67) );
  AND3X1 U363 ( .A(add_x_41_1_carry_12_), .B(cnt2[12]), .C(cnt2[13]), .Y(
        add_x_41_1_carry_14_) );
  AND2X1 U364 ( .A(add_x_41_1_carry_12_), .B(cnt2[12]), .Y(n387) );
  AOI2BB2X1 U365 ( .B0(n387), .B1(cnt2[13]), .A0N(n387), .A1N(cnt2[13]), .Y(
        N88) );
  NOR2BX1 U366 ( .AN(n99), .B(mode[0]), .Y(n103) );
  AOI2BB2X1 U367 ( .B0(cnt1[3]), .B1(add_x_41_0_carry_3_), .A0N(cnt1[3]), 
        .A1N(add_x_41_0_carry_3_), .Y(n388) );
  AO22X1 U368 ( .A0(cnt1[3]), .A1(n244), .B0(n388), .B1(n435), .Y(n349) );
  AND2X1 U369 ( .A(n392), .B(cnt1[19]), .Y(n389) );
  AOI2BB2X1 U370 ( .B0(n389), .B1(cnt1[20]), .A0N(n389), .A1N(cnt1[20]), .Y(
        n390) );
  AO22X1 U371 ( .A0(cnt1[20]), .A1(n244), .B0(n390), .B1(n435), .Y(n332) );
  INVX3 U373 ( .A(n394), .Y(add_x_41_1_carry_20_) );
  INVX1 U374 ( .A(n143), .Y(n93) );
  INVX1 U375 ( .A(n176), .Y(n92) );
  OR2X4 U376 ( .A(rst), .B(n98), .Y(n434) );
  ADDHX4 U377 ( .A(cnt2[1]), .B(cnt2[0]), .CO(add_x_41_1_carry_2_), .S(N76) );
  ADDHX4 U378 ( .A(cnt2[3]), .B(add_x_41_1_carry_3_), .CO(add_x_41_1_carry_4_), 
        .S(N78) );
  ADDHX4 U379 ( .A(cnt2[2]), .B(add_x_41_1_carry_2_), .CO(add_x_41_1_carry_3_), 
        .S(N77) );
  AOI2BB2X4 U380 ( .B0(add_x_41_1_carry_20_), .B1(cnt2[20]), .A0N(
        add_x_41_1_carry_20_), .A1N(cnt2[20]), .Y(N95) );
  XOR2XL U381 ( .A(cnt2[19]), .B(add_x_41_1_carry_19_), .Y(N94) );
  XOR2XL U382 ( .A(cnt2[12]), .B(add_x_41_1_carry_12_), .Y(N87) );
  ADDHX4 U383 ( .A(cnt2[14]), .B(add_x_41_1_carry_14_), .CO(
        add_x_41_1_carry_15_), .S(N89) );
  ADDHX4 U384 ( .A(cnt2[15]), .B(add_x_41_1_carry_15_), .CO(
        add_x_41_1_carry_16_), .S(N90) );
  AO22X4 U385 ( .A0(n44), .A1(N95), .B0(cnt2[20]), .B1(n245), .Y(n374) );
  NOR2X1 U386 ( .A(mode[2]), .B(n96), .Y(n99) );
  CLKINVX1 U387 ( .A(mode[0]), .Y(n97) );
  NOR3X1 U388 ( .A(n74), .B(n75), .C(n226), .Y(n231) );
  NAND2X1 U389 ( .A(n136), .B(n198), .Y(n226) );
  CLKINVX1 U390 ( .A(n148), .Y(n91) );
endmodule

